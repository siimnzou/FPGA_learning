module test
(
input a

output wire b
);

assign b =  a;

endmodule
