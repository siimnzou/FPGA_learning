/*********************************************************************
    字符信息获取模块，每个字符分别为128x128像素点
    通过之前模块传入的字符数（char_num）、字符x坐标、字符y坐标获取
    当前像素点的数据,传入pix_data模块，用于生成当前位置的rgb数据
**********************************************************************/
module CHAR_DATA
(
    input       clk,
    input       rst_n,
    input [9:0] char_x_loc,
    input [9:0] char_y_loc,
    input       char_data_req,
    input [3:0] char_num,

    output reg char_data 
);

reg [127:0] char [127:0] ;

// 不同数字取模 

always @(posedge clk or negedge rst_n) begin
    if (~rst_n)
        begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000000000000000000;
                char[22]   <=128'h0000000000001FFFFFF0000000000000;
                char[23]   <=128'h000000000001FFFFFFFF800000000000;
                char[24]   <=128'h00000000001FFFFFFFFFF80000000000;
                char[25]   <=128'h0000000000FFFFFFFFFFFE0000000000;
                char[26]   <=128'h0000000003FFFF00007FFFC000000000;
                char[27]   <=128'h000000000FFFF800000FFFF000000000;
                char[28]   <=128'h000000003FFFC0000001FFFC00000000;
                char[29]   <=128'h00000000FFFF800000007FFE00000000;
                char[30]   <=128'h00000001FFFE000000003FFF80000000;
                char[31]   <=128'h00000007FFFC000000001FFFE0000000;
                char[32]   <=128'h0000000FFFF00000000007FFF0000000;
                char[33]   <=128'h0000003FFFE00000000003FFF8000000;
                char[34]   <=128'h0000007FFFC00000000001FFFC000000;
                char[35]   <=128'h000000FFFF800000000001FFFE000000;
                char[36]   <=128'h000001FFFF000000000000FFFF000000;
                char[37]   <=128'h000003FFFE0000000000007FFF800000;
                char[38]   <=128'h000007FFFE0000000000003FFFC00000;
                char[39]   <=128'h000007FFFC0000000000003FFFE00000;
                char[40]   <=128'h00000FFFF80000000000001FFFF00000;
                char[41]   <=128'h00001FFFF80000000000001FFFF00000;
                char[42]   <=128'h00003FFFF00000000000000FFFF80000;
                char[43]   <=128'h00003FFFF00000000000000FFFFC0000;
                char[44]   <=128'h00007FFFE000000000000007FFFC0000;
                char[45]   <=128'h00007FFFE000000000000007FFFE0000;
                char[46]   <=128'h0000FFFFC000000000000007FFFE0000;
                char[47]   <=128'h0000FFFFC000000000000003FFFF0000;
                char[48]   <=128'h0001FFFF8000000000000003FFFF0000;
                char[49]   <=128'h0001FFFF8000000000000003FFFF0000;
                char[50]   <=128'h0003FFFF8000000000000003FFFF8000;
                char[51]   <=128'h0003FFFF8000000000000001FFFF8000;
                char[52]   <=128'h0003FFFF0000000000000001FFFF8000;
                char[53]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[54]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[55]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[56]   <=128'h0007FFFF0000000000000000FFFFC000;
                char[57]   <=128'h0007FFFE0000000000000000FFFFC000;
                char[58]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[59]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[60]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[61]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[62]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[63]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[64]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[65]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[66]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[67]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[68]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[69]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[70]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[71]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[72]   <=128'h0007FFFE0000000000000000FFFFC000;
                char[73]   <=128'h0007FFFF0000000000000000FFFFC000;
                char[74]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[75]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[76]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[77]   <=128'h0003FFFF0000000000000001FFFF8000;
                char[78]   <=128'h0003FFFF0000000000000001FFFF8000;
                char[79]   <=128'h0003FFFF8000000000000003FFFF8000;
                char[80]   <=128'h0003FFFF8000000000000003FFFF8000;
                char[81]   <=128'h0001FFFF8000000000000003FFFF0000;
                char[82]   <=128'h0001FFFFC000000000000003FFFF0000;
                char[83]   <=128'h0000FFFFC000000000000007FFFE0000;
                char[84]   <=128'h0000FFFFC000000000000007FFFE0000;
                char[85]   <=128'h00007FFFE000000000000007FFFC0000;
                char[86]   <=128'h00007FFFE00000000000000FFFFC0000;
                char[87]   <=128'h00003FFFF00000000000000FFFF80000;
                char[88]   <=128'h00003FFFF00000000000001FFFF80000;
                char[89]   <=128'h00001FFFF80000000000001FFFF00000;
                char[90]   <=128'h00000FFFF80000000000003FFFE00000;
                char[91]   <=128'h000007FFFC0000000000003FFFC00000;
                char[92]   <=128'h000003FFFE0000000000007FFF800000;
                char[93]   <=128'h000001FFFF000000000000FFFF800000;
                char[94]   <=128'h000000FFFF800000000001FFFF000000;
                char[95]   <=128'h0000007FFF800000000001FFFE000000;
                char[96]   <=128'h0000003FFFC00000000003FFF8000000;
                char[97]   <=128'h0000001FFFF00000000007FFF0000000;
                char[98]   <=128'h0000000FFFF8000000000FFFE0000000;
                char[99]   <=128'h00000003FFFC000000003FFF80000000;  
                char[100]  <=128'h00000001FFFF000000007FFF00000000;
                char[101]  <=128'h000000007FFF80000001FFFC00000000;
                char[102]  <=128'h000000001FFFE0000007FFF800000000;
                char[103]  <=128'h0000000007FFFC00003FFFE000000000;
                char[104]  <=128'h0000000001FFFFC003FFFF0000000000;
                char[105]  <=128'h00000000003FFFFFFFFFFC0000000000;
                char[106]  <=128'h000000000007FFFFFFFFE00000000000;
                char[107]  <=128'h0000000000007FFFFFFE000000000000;
                char[108]  <=128'h00000000000001FFFF80000000000000;
                char[109]  <=128'h00000000000000000000000000000000;
                char[110]  <=128'h00000000000000000000000000000000;
                char[111]  <=128'h00000000000000000000000000000000;
                char[112]  <=128'h00000000000000000000000000000000;
                char[113]  <=128'h00000000000000000000000000000000;
                char[114]  <=128'h00000000000000000000000000000000;
                char[115]  <=128'h00000000000000000000000000000000;
                char[116]  <=128'h00000000000000000000000000000000;
                char[117]  <=128'h00000000000000000000000000000000;
                char[118]  <=128'h00000000000000000000000000000000;
                char[119]  <=128'h00000000000000000000000000000000;
                char[120]  <=128'h00000000000000000000000000000000;
                char[121]  <=128'h00000000000000000000000000000000;
                char[122]  <=128'h00000000000000000000000000000000;
                char[123]  <=128'h00000000000000000000000000000000;
                char[124]  <=128'h00000000000000000000000000000000;
                char[125]  <=128'h00000000000000000000000000000000;
                char[126]  <=128'h00000000000000000000000000000000;
                char[127]  <=128'h00000000000000000000000000000000; 
        end
    else 
        case (char_num)
            4'd0:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000000000000000000;
                char[22]   <=128'h0000000000001FFFFFF0000000000000;
                char[23]   <=128'h000000000001FFFFFFFF800000000000;
                char[24]   <=128'h00000000001FFFFFFFFFF80000000000;
                char[25]   <=128'h0000000000FFFFFFFFFFFE0000000000;
                char[26]   <=128'h0000000003FFFF00007FFFC000000000;
                char[27]   <=128'h000000000FFFF800000FFFF000000000;
                char[28]   <=128'h000000003FFFC0000001FFFC00000000;
                char[29]   <=128'h00000000FFFF800000007FFE00000000;
                char[30]   <=128'h00000001FFFE000000003FFF80000000;
                char[31]   <=128'h00000007FFFC000000001FFFE0000000;
                char[32]   <=128'h0000000FFFF00000000007FFF0000000;
                char[33]   <=128'h0000003FFFE00000000003FFF8000000;
                char[34]   <=128'h0000007FFFC00000000001FFFC000000;
                char[35]   <=128'h000000FFFF800000000001FFFE000000;
                char[36]   <=128'h000001FFFF000000000000FFFF000000;
                char[37]   <=128'h000003FFFE0000000000007FFF800000;
                char[38]   <=128'h000007FFFE0000000000003FFFC00000;
                char[39]   <=128'h000007FFFC0000000000003FFFE00000;
                char[40]   <=128'h00000FFFF80000000000001FFFF00000;
                char[41]   <=128'h00001FFFF80000000000001FFFF00000;
                char[42]   <=128'h00003FFFF00000000000000FFFF80000;
                char[43]   <=128'h00003FFFF00000000000000FFFFC0000;
                char[44]   <=128'h00007FFFE000000000000007FFFC0000;
                char[45]   <=128'h00007FFFE000000000000007FFFE0000;
                char[46]   <=128'h0000FFFFC000000000000007FFFE0000;
                char[47]   <=128'h0000FFFFC000000000000003FFFF0000;
                char[48]   <=128'h0001FFFF8000000000000003FFFF0000;
                char[49]   <=128'h0001FFFF8000000000000003FFFF0000;
                char[50]   <=128'h0003FFFF8000000000000003FFFF8000;
                char[51]   <=128'h0003FFFF8000000000000001FFFF8000;
                char[52]   <=128'h0003FFFF0000000000000001FFFF8000;
                char[53]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[54]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[55]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[56]   <=128'h0007FFFF0000000000000000FFFFC000;
                char[57]   <=128'h0007FFFE0000000000000000FFFFC000;
                char[58]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[59]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[60]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[61]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[62]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[63]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[64]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[65]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[66]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[67]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[68]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[69]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[70]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[71]   <=128'h000FFFFE0000000000000000FFFFE000;
                char[72]   <=128'h0007FFFE0000000000000000FFFFC000;
                char[73]   <=128'h0007FFFF0000000000000000FFFFC000;
                char[74]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[75]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[76]   <=128'h0007FFFF0000000000000001FFFFC000;
                char[77]   <=128'h0003FFFF0000000000000001FFFF8000;
                char[78]   <=128'h0003FFFF0000000000000001FFFF8000;
                char[79]   <=128'h0003FFFF8000000000000003FFFF8000;
                char[80]   <=128'h0003FFFF8000000000000003FFFF8000;
                char[81]   <=128'h0001FFFF8000000000000003FFFF0000;
                char[82]   <=128'h0001FFFFC000000000000003FFFF0000;
                char[83]   <=128'h0000FFFFC000000000000007FFFE0000;
                char[84]   <=128'h0000FFFFC000000000000007FFFE0000;
                char[85]   <=128'h00007FFFE000000000000007FFFC0000;
                char[86]   <=128'h00007FFFE00000000000000FFFFC0000;
                char[87]   <=128'h00003FFFF00000000000000FFFF80000;
                char[88]   <=128'h00003FFFF00000000000001FFFF80000;
                char[89]   <=128'h00001FFFF80000000000001FFFF00000;
                char[90]   <=128'h00000FFFF80000000000003FFFE00000;
                char[91]   <=128'h000007FFFC0000000000003FFFC00000;
                char[92]   <=128'h000003FFFE0000000000007FFF800000;
                char[93]   <=128'h000001FFFF000000000000FFFF800000;
                char[94]   <=128'h000000FFFF800000000001FFFF000000;
                char[95]   <=128'h0000007FFF800000000001FFFE000000;
                char[96]   <=128'h0000003FFFC00000000003FFF8000000;
                char[97]   <=128'h0000001FFFF00000000007FFF0000000;
                char[98]   <=128'h0000000FFFF8000000000FFFE0000000;
                char[99]   <=128'h00000003FFFC000000003FFF80000000;  
                char[100]  <=128'h00000001FFFF000000007FFF00000000;
                char[101]  <=128'h000000007FFF80000001FFFC00000000;
                char[102]  <=128'h000000001FFFE0000007FFF800000000;
                char[103]  <=128'h0000000007FFFC00003FFFE000000000;
                char[104]  <=128'h0000000001FFFFC003FFFF0000000000;
                char[105]  <=128'h00000000003FFFFFFFFFFC0000000000;
                char[106]  <=128'h000000000007FFFFFFFFE00000000000;
                char[107]  <=128'h0000000000007FFFFFFE000000000000;
                char[108]  <=128'h00000000000001FFFF80000000000000;
                char[109]  <=128'h00000000000000000000000000000000;
                char[110]  <=128'h00000000000000000000000000000000;
                char[111]  <=128'h00000000000000000000000000000000;
                char[112]  <=128'h00000000000000000000000000000000;
                char[113]  <=128'h00000000000000000000000000000000;
                char[114]  <=128'h00000000000000000000000000000000;
                char[115]  <=128'h00000000000000000000000000000000;
                char[116]  <=128'h00000000000000000000000000000000;
                char[117]  <=128'h00000000000000000000000000000000;
                char[118]  <=128'h00000000000000000000000000000000;
                char[119]  <=128'h00000000000000000000000000000000;
                char[120]  <=128'h00000000000000000000000000000000;
                char[121]  <=128'h00000000000000000000000000000000;
                char[122]  <=128'h00000000000000000000000000000000;
                char[123]  <=128'h00000000000000000000000000000000;
                char[124]  <=128'h00000000000000000000000000000000;
                char[125]  <=128'h00000000000000000000000000000000;
                char[126]  <=128'h00000000000000000000000000000000;
                char[127]  <=128'h00000000000000000000000000000000; 
            end
        4'd1:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000F80000000000000;
                char[22]   <=128'h00000000000000001F80000000000000;
                char[23]   <=128'h00000000000000003F80000000000000;
                char[24]   <=128'h0000000000000000FF80000000000000;
                char[25]   <=128'h0000000000000003FF80000000000000;
                char[26]   <=128'h000000000000001FFF80000000000000;
                char[27]   <=128'h00000000000001FFFF80000000000000;
                char[28]   <=128'h0000000000007FFFFF80000000000000;
                char[29]   <=128'h00000007FFFFFFFFFF80000000000000;
                char[30]   <=128'h00000007FFFFFFFFFF80000000000000;
                char[31]   <=128'h00000007FFFFFFFFFF80000000000000;
                char[32]   <=128'h0000000000000FFFFF80000000000000;
                char[33]   <=128'h00000000000001FFFF80000000000000;
                char[34]   <=128'h00000000000000FFFF80000000000000;
                char[35]   <=128'h000000000000007FFF80000000000000;
                char[36]   <=128'h000000000000007FFF80000000000000;
                char[37]   <=128'h000000000000007FFF80000000000000;
                char[38]   <=128'h000000000000007FFF80000000000000;
                char[39]   <=128'h000000000000007FFF80000000000000;
                char[40]   <=128'h000000000000007FFF80000000000000;
                char[41]   <=128'h000000000000007FFF80000000000000;
                char[42]   <=128'h000000000000007FFF80000000000000;
                char[43]   <=128'h000000000000007FFF80000000000000;
                char[44]   <=128'h000000000000007FFF80000000000000;
                char[45]   <=128'h000000000000007FFF80000000000000;
                char[46]   <=128'h000000000000007FFF80000000000000;
                char[47]   <=128'h000000000000007FFF80000000000000;
                char[48]   <=128'h000000000000007FFF80000000000000;
                char[49]   <=128'h000000000000007FFF80000000000000;
                char[50]   <=128'h000000000000007FFF80000000000000;
                char[51]   <=128'h000000000000007FFF80000000000000;
                char[52]   <=128'h000000000000007FFF80000000000000;
                char[53]   <=128'h000000000000007FFF80000000000000;
                char[54]   <=128'h000000000000007FFF80000000000000;
                char[55]   <=128'h000000000000007FFF80000000000000;
                char[56]   <=128'h000000000000007FFF80000000000000;
                char[57]   <=128'h000000000000007FFF80000000000000;
                char[58]   <=128'h000000000000007FFF80000000000000;
                char[59]   <=128'h000000000000007FFF80000000000000;
                char[60]   <=128'h000000000000007FFF80000000000000;
                char[61]   <=128'h000000000000007FFF80000000000000;
                char[62]   <=128'h000000000000007FFF80000000000000;
                char[63]   <=128'h000000000000007FFF80000000000000;
                char[64]   <=128'h000000000000007FFF80000000000000;
                char[65]   <=128'h000000000000007FFF80000000000000;
                char[66]   <=128'h000000000000007FFF80000000000000;
                char[67]   <=128'h000000000000007FFF80000000000000;
                char[68]   <=128'h000000000000007FFF80000000000000;
                char[69]   <=128'h000000000000007FFF80000000000000;
                char[70]   <=128'h000000000000007FFF80000000000000;
                char[71]   <=128'h000000000000007FFF80000000000000;
                char[72]   <=128'h000000000000007FFF80000000000000;
                char[73]   <=128'h000000000000007FFF80000000000000;
                char[74]   <=128'h000000000000007FFF80000000000000;
                char[75]   <=128'h000000000000007FFF80000000000000;
                char[76]   <=128'h000000000000007FFF80000000000000;
                char[77]   <=128'h000000000000007FFF80000000000000;
                char[78]   <=128'h000000000000007FFF80000000000000;
                char[79]   <=128'h000000000000007FFF80000000000000;
                char[80]   <=128'h000000000000007FFF80000000000000;
                char[81]   <=128'h000000000000007FFF80000000000000;
                char[82]   <=128'h000000000000007FFF80000000000000;
                char[83]   <=128'h000000000000007FFF80000000000000;
                char[84]   <=128'h000000000000007FFF80000000000000;
                char[85]   <=128'h000000000000007FFF80000000000000;
                char[86]   <=128'h000000000000007FFF80000000000000;
                char[87]   <=128'h000000000000007FFF80000000000000;
                char[88]   <=128'h000000000000007FFF80000000000000;
                char[89]   <=128'h000000000000007FFF80000000000000;
                char[90]   <=128'h000000000000007FFF80000000000000;
                char[91]   <=128'h000000000000007FFF80000000000000;
                char[92]   <=128'h000000000000007FFF80000000000000;
                char[93]   <=128'h000000000000007FFF80000000000000;
                char[94]   <=128'h000000000000007FFF80000000000000;
                char[95]   <=128'h000000000000007FFF80000000000000;
                char[96]   <=128'h000000000000007FFF80000000000000;
                char[97]   <=128'h000000000000007FFF80000000000000;
                char[98]   <=128'h000000000000007FFF80000000000000;
                char[99]   <=128'h00000000000000FFFFC0000000000000;   
                char[100]  <=128'h00000000000000FFFFC0000000000000; 
                char[101]  <=128'h00000000000001FFFFE0000000000000; 
                char[102]  <=128'h00000000000007FFFFF8000000000000; 
                char[103]  <=128'h0000000000001FFFFFFE000000000000; 
                char[104]  <=128'h000000000001FFFFFFFFF00000000000; 
                char[105]  <=128'h00000007FFFFFFFFFFFFFFFFFC000000; 
                char[106]  <=128'h00000007FFFFFFFFFFFFFFFFFC000000; 
                char[107]  <=128'h00000007FFFFFFFFFFFFFFFFFC000000; 
                char[108]  <=128'h00000000000000000000000000000000; 
                char[109]  <=128'h00000000000000000000000000000000; 
                char[110]  <=128'h00000000000000000000000000000000; 
                char[111]  <=128'h00000000000000000000000000000000; 
                char[112]  <=128'h00000000000000000000000000000000; 
                char[113]  <=128'h00000000000000000000000000000000; 
                char[114]  <=128'h00000000000000000000000000000000; 
                char[115]  <=128'h00000000000000000000000000000000; 
                char[116]  <=128'h00000000000000000000000000000000; 
                char[117]  <=128'h00000000000000000000000000000000; 
                char[118]  <=128'h00000000000000000000000000000000; 
                char[119]  <=128'h00000000000000000000000000000000; 
                char[120]  <=128'h00000000000000000000000000000000; 
                char[121]  <=128'h00000000000000000000000000000000; 
                char[122]  <=128'h00000000000000000000000000000000; 
                char[123]  <=128'h00000000000000000000000000000000; 
                char[124]  <=128'h00000000000000000000000000000000; 
                char[125]  <=128'h00000000000000000000000000000000; 
                char[126]  <=128'h00000000000000000000000000000000; 
                char[127]  <=128'h00000000000000000000000000000000;  
            end
            4'd2:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000000000000000000;
                char[22]   <=128'h0000000000007FFFFFFF800000000000;
                char[23]   <=128'h00000000001FFFFFFFFFFE0000000000;
                char[24]   <=128'h0000000001FFFFFFFFFFFFE000000000;
                char[25]   <=128'h000000001FFFF00001FFFFFC00000000;
                char[26]   <=128'h00000000FFFC0000000FFFFF00000000;
                char[27]   <=128'h00000003FFE000000000FFFFE0000000;
                char[28]   <=128'h0000001FFF00000000001FFFF0000000;
                char[29]   <=128'h0000007FFC000000000007FFFC000000;
                char[30]   <=128'h000000FFF0000000000003FFFE000000;
                char[31]   <=128'h000003FFE0000000000000FFFF800000;
                char[32]   <=128'h000007FFC00000000000007FFFC00000;
                char[33]   <=128'h00000FFF800000000000003FFFE00000;
                char[34]   <=128'h00001FFF000000000000003FFFE00000;
                char[35]   <=128'h00003FFF000000000000001FFFF00000;
                char[36]   <=128'h00003FFF000000000000001FFFF80000;
                char[37]   <=128'h00007FFF000000000000000FFFF80000;
                char[38]   <=128'h00007FFF800000000000000FFFF80000;
                char[39]   <=128'h0000FFFF8000000000000007FFFC0000;
                char[40]   <=128'h0000FFFFC000000000000007FFFC0000;
                char[41]   <=128'h0000FFFFF000000000000007FFFC0000;
                char[42]   <=128'h0000FFFFF800000000000007FFFC0000;
                char[43]   <=128'h0000FFFFFC00000000000007FFFC0000;
                char[44]   <=128'h0000FFFFFE00000000000007FFFC0000;
                char[45]   <=128'h0000FFFFFE00000000000007FFFC0000;
                char[46]   <=128'h00007FFFFE00000000000007FFF80000;
                char[47]   <=128'h00003FFFFC0000000000000FFFF80000;
                char[48]   <=128'h00001FFFFC0000000000000FFFF80000;
                char[49]   <=128'h000007FFF00000000000001FFFF00000;
                char[50]   <=128'h00000000000000000000001FFFF00000;
                char[51]   <=128'h00000000000000000000003FFFE00000;
                char[52]   <=128'h00000000000000000000003FFFC00000;
                char[53]   <=128'h00000000000000000000007FFF800000;
                char[54]   <=128'h0000000000000000000000FFFF800000;
                char[55]   <=128'h0000000000000000000001FFFF000000;
                char[56]   <=128'h0000000000000000000003FFFC000000;
                char[57]   <=128'h0000000000000000000007FFF8000000;
                char[58]   <=128'h000000000000000000000FFFF0000000;
                char[59]   <=128'h000000000000000000001FFFE0000000;
                char[60]   <=128'h000000000000000000007FFF80000000;
                char[61]   <=128'h00000000000000000000FFFF00000000;
                char[62]   <=128'h00000000000000000001FFFC00000000;
                char[63]   <=128'h00000000000000000007FFF000000000;
                char[64]   <=128'h0000000000000000000FFFC000000000;
                char[65]   <=128'h0000000000000000003FFF0000000000;
                char[66]   <=128'h0000000000000000007FFC0000000000;
                char[67]   <=128'h000000000000000001FFF00000000000;
                char[68]   <=128'h000000000000000007FFC00000000000;
                char[69]   <=128'h00000000000000000FFF000000000000;
                char[70]   <=128'h00000000000000003FFC000000000000;
                char[71]   <=128'h0000000000000000FFF0000000000000;
                char[72]   <=128'h0000000000000003FFC0000000000000;
                char[73]   <=128'h000000000000000FFF00000000000000;
                char[74]   <=128'h000000000000003FFC00000000000000;
                char[75]   <=128'h00000000000000FFF000000000000000;
                char[76]   <=128'h00000000000003FFC000000000000000;
                char[77]   <=128'h0000000000000FFF0000000000000000;
                char[78]   <=128'h0000000000003FFC0000000000000000;
                char[79]   <=128'h000000000000FFF00000000000000000;
                char[80]   <=128'h000000000003FFC00000000000000000;
                char[81]   <=128'h000000000007FF000000000000000000;
                char[82]   <=128'h00000000001FFC000000000000000000;
                char[83]   <=128'h00000000007FF0000000000000000000;
                char[84]   <=128'h0000000001FFC0000000000000000000;
                char[85]   <=128'h0000000007FF00000000000000000000;
                char[86]   <=128'h000000001FFE000000000000003F0000;
                char[87]   <=128'h000000003FF8000000000000003F0000;
                char[88]   <=128'h00000000FFE0000000000000007E0000;
                char[89]   <=128'h00000003FF80000000000000007E0000;
                char[90]   <=128'h00000007FE0000000000000000FE0000;
                char[91]   <=128'h0000001FFC0000000000000000FE0000;
                char[92]   <=128'h0000007FF00000000000000001FC0000;
                char[93]   <=128'h000000FFC00000000000000003FC0000;
                char[94]   <=128'h000003FF800000000000000007FC0000;
                char[95]   <=128'h000007FE00000000000000000FF80000;
                char[96]   <=128'h00001FF800000000000000001FF80000;
                char[97]   <=128'h00003FF000000000000000007FF80000;
                char[98]   <=128'h00007FC00000000000000001FFF80000;
                char[99]   <=128'h0001FF80000000000000000FFFF00000;   
                char[100]  <=128'h0003FFFFFFFFFFFFFFFFFFFFFFF00000; 
                char[101]  <=128'h0007FFFFFFFFFFFFFFFFFFFFFFF00000; 
                char[102]  <=128'h0007FFFFFFFFFFFFFFFFFFFFFFF00000; 
                char[103]  <=128'h0007FFFFFFFFFFFFFFFFFFFFFFE00000; 
                char[104]  <=128'h0007FFFFFFFFFFFFFFFFFFFFFFE00000; 
                char[105]  <=128'h0007FFFFFFFFFFFFFFFFFFFFFFE00000; 
                char[106]  <=128'h0007FFFFFFFFFFFFFFFFFFFFFFC00000; 
                char[107]  <=128'h0007FFFFFFFFFFFFFFFFFFFFFFC00000; 
                char[108]  <=128'h00000000000000000000000000000000; 
                char[109]  <=128'h00000000000000000000000000000000; 
                char[110]  <=128'h00000000000000000000000000000000; 
                char[111]  <=128'h00000000000000000000000000000000; 
                char[112]  <=128'h00000000000000000000000000000000; 
                char[113]  <=128'h00000000000000000000000000000000; 
                char[114]  <=128'h00000000000000000000000000000000; 
                char[115]  <=128'h00000000000000000000000000000000; 
                char[116]  <=128'h00000000000000000000000000000000; 
                char[117]  <=128'h00000000000000000000000000000000; 
                char[118]  <=128'h00000000000000000000000000000000; 
                char[119]  <=128'h00000000000000000000000000000000; 
                char[120]  <=128'h00000000000000000000000000000000; 
                char[121]  <=128'h00000000000000000000000000000000; 
                char[122]  <=128'h00000000000000000000000000000000; 
                char[123]  <=128'h00000000000000000000000000000000; 
                char[124]  <=128'h00000000000000000000000000000000; 
                char[125]  <=128'h00000000000000000000000000000000; 
                char[126]  <=128'h00000000000000000000000000000000; 
                char[127]  <=128'h00000000000000000000000000000000; 
            end 
            4'd3:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000000000000000000;
                char[22]   <=128'h000000000003FFFFFFF0000000000000;
                char[23]   <=128'h00000000007FFFFFFFFF800000000000;
                char[24]   <=128'h0000000007FFFFFFFFFFF80000000000;
                char[25]   <=128'h000000007FFF80003FFFFF0000000000;
                char[26]   <=128'h00000003FFE0000000FFFFC000000000;
                char[27]   <=128'h0000000FFE000000001FFFF800000000;
                char[28]   <=128'h0000003FF80000000007FFFC00000000;
                char[29]   <=128'h000000FFE00000000001FFFF00000000;
                char[30]   <=128'h000001FFE000000000007FFFC0000000;
                char[31]   <=128'h000007FFC000000000003FFFE0000000;
                char[32]   <=128'h00000FFFC000000000001FFFF0000000;
                char[33]   <=128'h00000FFFC000000000000FFFF8000000;
                char[34]   <=128'h00001FFFC0000000000007FFFC000000;
                char[35]   <=128'h00001FFFC0000000000003FFFE000000;
                char[36]   <=128'h00003FFFE0000000000003FFFF000000;
                char[37]   <=128'h00003FFFF0000000000001FFFF000000;
                char[38]   <=128'h00003FFFF8000000000001FFFF800000;
                char[39]   <=128'h00003FFFFC000000000000FFFF800000;
                char[40]   <=128'h00003FFFFC000000000000FFFF800000;
                char[41]   <=128'h00001FFFFC000000000000FFFF800000;
                char[42]   <=128'h00001FFFF8000000000000FFFF800000;
                char[43]   <=128'h000007FFF8000000000000FFFF800000;
                char[44]   <=128'h000001FFE0000000000000FFFF800000;
                char[45]   <=128'h0000000000000000000000FFFF000000;
                char[46]   <=128'h0000000000000000000001FFFF000000;
                char[47]   <=128'h0000000000000000000001FFFE000000;
                char[48]   <=128'h0000000000000000000001FFFE000000;
                char[49]   <=128'h0000000000000000000003FFFC000000;
                char[50]   <=128'h0000000000000000000007FFF8000000;
                char[51]   <=128'h000000000000000000000FFFF0000000;
                char[52]   <=128'h000000000000000000001FFFE0000000;
                char[53]   <=128'h000000000000000000003FFFC0000000;
                char[54]   <=128'h000000000000000000007FFF00000000;
                char[55]   <=128'h00000000000000000001FFFE00000000;
                char[56]   <=128'h00000000000000000007FFF800000000;
                char[57]   <=128'h0000000000000000003FFFC000000000;
                char[58]   <=128'h000000000000000001FFFE0000000000;
                char[59]   <=128'h00000000000000007FFFF00000000000;
                char[60]   <=128'h0000000000007FFFFFFF000000000000;
                char[61]   <=128'h0000000000007FFFFFC0000000000000;
                char[62]   <=128'h0000000000007FFFFFFE000000000000;
                char[63]   <=128'h0000000000007FFFFFFFE00000000000;
                char[64]   <=128'h0000000000000001FFFFFE0000000000;
                char[65]   <=128'h000000000000000000FFFFE000000000;
                char[66]   <=128'h00000000000000000007FFFC00000000;
                char[67]   <=128'h00000000000000000000FFFF00000000;
                char[68]   <=128'h000000000000000000001FFFC0000000;
                char[69]   <=128'h000000000000000000000FFFF0000000;
                char[70]   <=128'h0000000000000000000003FFFC000000;
                char[71]   <=128'h0000000000000000000001FFFE000000;
                char[72]   <=128'h00000000000000000000007FFF800000;
                char[73]   <=128'h00000000000000000000003FFFC00000;
                char[74]   <=128'h00000000000000000000001FFFE00000;
                char[75]   <=128'h00000000000000000000001FFFF00000;
                char[76]   <=128'h00000000000000000000000FFFF80000;
                char[77]   <=128'h000000000000000000000007FFF80000;
                char[78]   <=128'h000000000000000000000007FFFC0000;
                char[79]   <=128'h000000000000000000000007FFFE0000;
                char[80]   <=128'h000000000000000000000003FFFE0000;
                char[81]   <=128'h000000000000000000000003FFFE0000;
                char[82]   <=128'h000000000000000000000003FFFF0000;
                char[83]   <=128'h000000000000000000000003FFFF0000;
                char[84]   <=128'h000000000000000000000003FFFF0000;
                char[85]   <=128'h000001FF0000000000000003FFFF0000;
                char[86]   <=128'h00000FFFC000000000000003FFFF0000;
                char[87]   <=128'h00001FFFF000000000000003FFFF0000;
                char[88]   <=128'h00007FFFF800000000000003FFFF0000;
                char[89]   <=128'h0000FFFFF800000000000007FFFE0000;
                char[90]   <=128'h0001FFFFFC00000000000007FFFE0000;
                char[91]   <=128'h0001FFFFFC00000000000007FFFC0000;
                char[92]   <=128'h0001FFFFFC0000000000000FFFFC0000;
                char[93]   <=128'h0001FFFFF80000000000000FFFF80000;
                char[94]   <=128'h0001FFFFF80000000000001FFFF00000;
                char[95]   <=128'h0000FFFFF00000000000003FFFE00000;
                char[96]   <=128'h0000FFFFE00000000000003FFFC00000;
                char[97]   <=128'h00007FFFC00000000000007FFF800000;
                char[98]   <=128'h00003FFFC0000000000000FFFE000000;
                char[99]   <=128'h00001FFFC0000000000003FFFC000000;   
                char[100]  <=128'h000007FFE0000000000007FFF0000000; 
                char[101]  <=128'h000003FFF000000000001FFFC0000000; 
                char[102]  <=128'h000000FFFC0000000000FFFF00000000; 
                char[103]  <=128'h0000001FFFC000000007FFFC00000000; 
                char[104]  <=128'h00000007FFFC000000FFFFF000000000; 
                char[105]  <=128'h00000000FFFFFFFFFFFFFF0000000000; 
                char[106]  <=128'h000000000FFFFFFFFFFFF80000000000; 
                char[107]  <=128'h00000000007FFFFFFFFE000000000000; 
                char[108]  <=128'h000000000000FFFFFE00000000000000; 
                char[109]  <=128'h00000000000000000000000000000000; 
                char[110]  <=128'h00000000000000000000000000000000; 
                char[111]  <=128'h00000000000000000000000000000000; 
                char[112]  <=128'h00000000000000000000000000000000; 
                char[113]  <=128'h00000000000000000000000000000000; 
                char[114]  <=128'h00000000000000000000000000000000; 
                char[115]  <=128'h00000000000000000000000000000000; 
                char[116]  <=128'h00000000000000000000000000000000; 
                char[117]  <=128'h00000000000000000000000000000000; 
                char[118]  <=128'h00000000000000000000000000000000; 
                char[119]  <=128'h00000000000000000000000000000000; 
                char[120]  <=128'h00000000000000000000000000000000; 
                char[121]  <=128'h00000000000000000000000000000000; 
                char[122]  <=128'h00000000000000000000000000000000; 
                char[123]  <=128'h00000000000000000000000000000000; 
                char[124]  <=128'h00000000000000000000000000000000; 
                char[125]  <=128'h00000000000000000000000000000000; 
                char[126]  <=128'h00000000000000000000000000000000; 
                char[127]  <=128'h00000000000000000000000000000000;  
            end
            4'd4:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h000000000000000000003FF000000000;
                char[22]   <=128'h000000000000000000007FF000000000;
                char[23]   <=128'h00000000000000000001FFF000000000;
                char[24]   <=128'h00000000000000000003FFF000000000;
                char[25]   <=128'h00000000000000000007FFF000000000;
                char[26]   <=128'h0000000000000000000FFFF000000000;
                char[27]   <=128'h0000000000000000003FFFF000000000;
                char[28]   <=128'h0000000000000000007FFFF000000000;
                char[29]   <=128'h000000000000000000FFFFF000000000;
                char[30]   <=128'h000000000000000001FFFFF000000000;
                char[31]   <=128'h000000000000000007FFFFF000000000;
                char[32]   <=128'h00000000000000000FFFFFF000000000;
                char[33]   <=128'h00000000000000001FFFFFF000000000;
                char[34]   <=128'h00000000000000003FCFFFF000000000;
                char[35]   <=128'h0000000000000000FF8FFFF000000000;
                char[36]   <=128'h0000000000000001FF0FFFF000000000;
                char[37]   <=128'h0000000000000003FE0FFFF000000000;
                char[38]   <=128'h0000000000000007F80FFFF000000000;
                char[39]   <=128'h000000000000001FF00FFFF000000000;
                char[40]   <=128'h000000000000003FE00FFFF000000000;
                char[41]   <=128'h000000000000007FC00FFFF000000000;
                char[42]   <=128'h00000000000000FF000FFFF000000000;
                char[43]   <=128'h00000000000003FE000FFFF000000000;
                char[44]   <=128'h00000000000007FC000FFFF000000000;
                char[45]   <=128'h0000000000000FF0000FFFF000000000;
                char[46]   <=128'h0000000000001FE0000FFFF000000000;
                char[47]   <=128'h0000000000007FC0000FFFF000000000;
                char[48]   <=128'h000000000000FF80000FFFF000000000;
                char[49]   <=128'h000000000001FE00000FFFF000000000;
                char[50]   <=128'h000000000007FC00000FFFF000000000;
                char[51]   <=128'h00000000000FF800000FFFF000000000;
                char[52]   <=128'h00000000001FF000000FFFF000000000;
                char[53]   <=128'h00000000003FC000000FFFF000000000;
                char[54]   <=128'h0000000000FF8000000FFFF000000000;
                char[55]   <=128'h0000000001FF0000000FFFF000000000;
                char[56]   <=128'h0000000003FE0000000FFFF000000000;
                char[57]   <=128'h0000000007F80000000FFFF000000000;
                char[58]   <=128'h000000001FF00000000FFFF000000000;
                char[59]   <=128'h000000003FE00000000FFFF000000000;
                char[60]   <=128'h000000007F800000000FFFF000000000;
                char[61]   <=128'h00000000FF000000000FFFF000000000;
                char[62]   <=128'h00000003FE000000000FFFF000000000;
                char[63]   <=128'h00000007FC000000000FFFF000000000;
                char[64]   <=128'h0000000FF0000000000FFFF000000000;
                char[65]   <=128'h0000001FE0000000000FFFF000000000;
                char[66]   <=128'h0000007FC0000000000FFFF000000000;
                char[67]   <=128'h000000FF80000000000FFFF000000000;
                char[68]   <=128'h000001FE00000000000FFFF000000000;
                char[69]   <=128'h000003FC00000000000FFFF000000000;
                char[70]   <=128'h00000FF800000000000FFFF000000000;
                char[71]   <=128'h00001FF000000000000FFFF000000000;
                char[72]   <=128'h00003FC000000000000FFFF000000000;
                char[73]   <=128'h00007F8000000000000FFFF000000000;
                char[74]   <=128'h0001FF0000000000000FFFF000000000;
                char[75]   <=128'h0003FC0000000000000FFFF000000000;
                char[76]   <=128'h0007F80000000000000FFFF000000000;
                char[77]   <=128'h000FF00000000000000FFFF000000000;
                char[78]   <=128'h003FE00000000000000FFFF000000000;
                char[79]   <=128'h007FFFFFFFFFFFFFFFFFFFFFFFFFFE00;
                char[80]   <=128'h007FFFFFFFFFFFFFFFFFFFFFFFFFFE00;
                char[81]   <=128'h007FFFFFFFFFFFFFFFFFFFFFFFFFFE00;
                char[82]   <=128'h0000000000000000000FFFF000000000;
                char[83]   <=128'h0000000000000000000FFFF000000000;
                char[84]   <=128'h0000000000000000000FFFF000000000;
                char[85]   <=128'h0000000000000000000FFFF000000000;
                char[86]   <=128'h0000000000000000000FFFF000000000;
                char[87]   <=128'h0000000000000000000FFFF000000000;
                char[88]   <=128'h0000000000000000000FFFF000000000;
                char[89]   <=128'h0000000000000000000FFFF000000000;
                char[90]   <=128'h0000000000000000000FFFF000000000;
                char[91]   <=128'h0000000000000000000FFFF000000000;
                char[92]   <=128'h0000000000000000000FFFF000000000;
                char[93]   <=128'h0000000000000000000FFFF000000000;
                char[94]   <=128'h0000000000000000000FFFF000000000;
                char[95]   <=128'h0000000000000000000FFFF000000000;
                char[96]   <=128'h0000000000000000000FFFF000000000;
                char[97]   <=128'h0000000000000000000FFFF000000000;
                char[98]   <=128'h0000000000000000000FFFF000000000;
                char[99]   <=128'h0000000000000000000FFFF000000000;   
                char[100]  <=128'h0000000000000000000FFFF000000000; 
                char[101]  <=128'h0000000000000000001FFFF800000000; 
                char[102]  <=128'h0000000000000000003FFFFC00000000; 
                char[103]  <=128'h000000000000000000FFFFFF00000000; 
                char[104]  <=128'h000000000000000007FFFFFFF0000000; 
                char[105]  <=128'h0000000000003FFFFFFFFFFFFFFFF000; 
                char[106]  <=128'h0000000000003FFFFFFFFFFFFFFFF000; 
                char[107]  <=128'h0000000000003FFFFFFFFFFFFFFFF000; 
                char[108]  <=128'h00000000000000000000000000000000; 
                char[109]  <=128'h00000000000000000000000000000000; 
                char[110]  <=128'h00000000000000000000000000000000; 
                char[111]  <=128'h00000000000000000000000000000000; 
                char[112]  <=128'h00000000000000000000000000000000; 
                char[113]  <=128'h00000000000000000000000000000000; 
                char[114]  <=128'h00000000000000000000000000000000; 
                char[115]  <=128'h00000000000000000000000000000000; 
                char[116]  <=128'h00000000000000000000000000000000; 
                char[117]  <=128'h00000000000000000000000000000000; 
                char[118]  <=128'h00000000000000000000000000000000; 
                char[119]  <=128'h00000000000000000000000000000000; 
                char[120]  <=128'h00000000000000000000000000000000; 
                char[121]  <=128'h00000000000000000000000000000000; 
                char[122]  <=128'h00000000000000000000000000000000; 
                char[123]  <=128'h00000000000000000000000000000000; 
                char[124]  <=128'h00000000000000000000000000000000; 
                char[125]  <=128'h00000000000000000000000000000000; 
                char[126]  <=128'h00000000000000000000000000000000; 
                char[127]  <=128'h00000000000000000000000000000000;  
            end
            4'd5:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000000000000000000;
                char[22]   <=128'h0000001FFFFFFFFFFFFFFFFFFFF80000;
                char[23]   <=128'h0000001FFFFFFFFFFFFFFFFFFFF80000;
                char[24]   <=128'h0000001FFFFFFFFFFFFFFFFFFFF00000;
                char[25]   <=128'h0000001FFFFFFFFFFFFFFFFFFFF00000;
                char[26]   <=128'h0000001FFFFFFFFFFFFFFFFFFFE00000;
                char[27]   <=128'h0000003FFFFFFFFFFFFFFFFFFFE00000;
                char[28]   <=128'h0000003FFFFFFFFFFFFFFFFFFFE00000;
                char[29]   <=128'h0000003FFFFFFFFFFFFFFFFFFFC00000;
                char[30]   <=128'h0000003FC00000000000000000000000;
                char[31]   <=128'h0000003FC00000000000000000000000;
                char[32]   <=128'h0000003FC00000000000000000000000;
                char[33]   <=128'h0000003FC00000000000000000000000;
                char[34]   <=128'h0000003F800000000000000000000000;
                char[35]   <=128'h0000003F800000000000000000000000;
                char[36]   <=128'h0000007F800000000000000000000000;
                char[37]   <=128'h0000007F800000000000000000000000;
                char[38]   <=128'h0000007F800000000000000000000000;
                char[39]   <=128'h0000007F800000000000000000000000;
                char[40]   <=128'h0000007F800000000000000000000000;
                char[41]   <=128'h0000007F800000000000000000000000;
                char[42]   <=128'h0000007F000000000000000000000000;
                char[43]   <=128'h0000007F000000000000000000000000;
                char[44]   <=128'h0000007F000000000000000000000000;
                char[45]   <=128'h000000FF000000000000000000000000;
                char[46]   <=128'h000000FF000000000000000000000000;
                char[47]   <=128'h000000FF000000000000000000000000;
                char[48]   <=128'h000000FF000000000000000000000000;
                char[49]   <=128'h000000FF000000000000000000000000;
                char[50]   <=128'h000000FF000000000000000000000000;
                char[51]   <=128'h000000FE000000000000000000000000;
                char[52]   <=128'h000000FE000000000000000000000000;
                char[53]   <=128'h000000FE0000003FFFFC000000000000;
                char[54]   <=128'h000001FE00007FFFFFFFF80000000000;
                char[55]   <=128'h000001FE0007FFFFFFFFFF8000000000;
                char[56]   <=128'h000001FE003FFFFFFFFFFFF000000000;
                char[57]   <=128'h000001FE00FFFFFFFFFFFFFE00000000;
                char[58]   <=128'h000001FE07FFFE00007FFFFF80000000;
                char[59]   <=128'h000001FC0FFF00000003FFFFE0000000;
                char[60]   <=128'h000001FC3FF0000000007FFFF0000000;
                char[61]   <=128'h000001FCFFC0000000001FFFFC000000;
                char[62]   <=128'h000001FDFE000000000007FFFE000000;
                char[63]   <=128'h000003FFFC000000000001FFFF800000;
                char[64]   <=128'h000003FFF0000000000000FFFFC00000;
                char[65]   <=128'h000003FFE00000000000007FFFE00000;
                char[66]   <=128'h000003FF800000000000003FFFE00000;
                char[67]   <=128'h000003FF000000000000001FFFF00000;
                char[68]   <=128'h00000000000000000000001FFFF80000;
                char[69]   <=128'h00000000000000000000000FFFF80000;
                char[70]   <=128'h000000000000000000000007FFFC0000;
                char[71]   <=128'h000000000000000000000007FFFC0000;
                char[72]   <=128'h000000000000000000000003FFFE0000;
                char[73]   <=128'h000000000000000000000003FFFE0000;
                char[74]   <=128'h000000000000000000000003FFFE0000;
                char[75]   <=128'h000000000000000000000003FFFF0000;
                char[76]   <=128'h000000000000000000000001FFFF0000;
                char[77]   <=128'h000000000000000000000001FFFF0000;
                char[78]   <=128'h000000000000000000000001FFFF0000;
                char[79]   <=128'h000000000000000000000001FFFF0000;
                char[80]   <=128'h000000000000000000000001FFFF0000;
                char[81]   <=128'h000000000000000000000001FFFF0000;
                char[82]   <=128'h000000000000000000000001FFFF0000;
                char[83]   <=128'h000000000000000000000001FFFF0000;
                char[84]   <=128'h000007FFC000000000000001FFFF0000;
                char[85]   <=128'h00001FFFF000000000000001FFFE0000;
                char[86]   <=128'h00007FFFF800000000000003FFFE0000;
                char[87]   <=128'h0000FFFFFC00000000000003FFFE0000;
                char[88]   <=128'h0000FFFFFC00000000000003FFFC0000;
                char[89]   <=128'h0001FFFFFC00000000000003FFFC0000;
                char[90]   <=128'h0001FFFFFC00000000000007FFF80000;
                char[91]   <=128'h0001FFFFF800000000000007FFF80000;
                char[92]   <=128'h0001FFFFF00000000000000FFFF00000;
                char[93]   <=128'h0001FFFFE00000000000000FFFF00000;
                char[94]   <=128'h0000FFFFC00000000000001FFFE00000;
                char[95]   <=128'h0000FFFF800000000000003FFFC00000;
                char[96]   <=128'h00007FFF000000000000007FFF800000;
                char[97]   <=128'h00003FFF00000000000000FFFF000000;
                char[98]   <=128'h00001FFF00000000000001FFFE000000;
                char[99]   <=128'h00000FFF80000000000003FFFC000000;   
                char[100]  <=128'h000003FFC000000000000FFFF0000000; 
                char[101]  <=128'h000000FFE000000000003FFFE0000000; 
                char[102]  <=128'h0000003FFC0000000000FFFF80000000; 
                char[103]  <=128'h0000000FFFC000000007FFFE00000000; 
                char[104]  <=128'h00000001FFFE0000007FFFF000000000; 
                char[105]  <=128'h000000003FFFFFFFFFFFFF8000000000; 
                char[106]  <=128'h0000000003FFFFFFFFFFFC0000000000; 
                char[107]  <=128'h00000000001FFFFFFFFF800000000000; 
                char[108]  <=128'h0000000000003FFFFF80000000000000; 
                char[109]  <=128'h00000000000000000000000000000000; 
                char[110]  <=128'h00000000000000000000000000000000; 
                char[111]  <=128'h00000000000000000000000000000000; 
                char[112]  <=128'h00000000000000000000000000000000; 
                char[113]  <=128'h00000000000000000000000000000000; 
                char[114]  <=128'h00000000000000000000000000000000; 
                char[115]  <=128'h00000000000000000000000000000000; 
                char[116]  <=128'h00000000000000000000000000000000; 
                char[117]  <=128'h00000000000000000000000000000000; 
                char[118]  <=128'h00000000000000000000000000000000; 
                char[119]  <=128'h00000000000000000000000000000000; 
                char[120]  <=128'h00000000000000000000000000000000; 
                char[121]  <=128'h00000000000000000000000000000000; 
                char[122]  <=128'h00000000000000000000000000000000; 
                char[123]  <=128'h00000000000000000000000000000000; 
                char[124]  <=128'h00000000000000000000000000000000; 
                char[125]  <=128'h00000000000000000000000000000000; 
                char[126]  <=128'h00000000000000000000000000000000; 
                char[127]  <=128'h00000000000000000000000000000000;  
            end
            4'd6:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000000000000000000;
                char[22]   <=128'h000000000000001FFFFFFF0000000000;
                char[23]   <=128'h00000000000003FFFFFFFFF000000000;
                char[24]   <=128'h0000000000007FFFFFFFFFFE00000000;
                char[25]   <=128'h000000000003FFFF0000FFFFC0000000;
                char[26]   <=128'h00000000001FFFC000000FFFF0000000;
                char[27]   <=128'h0000000000FFFC00000007FFF8000000;
                char[28]   <=128'h0000000003FFE000000003FFFE000000;
                char[29]   <=128'h000000000FFF8000000003FFFF000000;
                char[30]   <=128'h000000003FFE0000000003FFFF800000;
                char[31]   <=128'h00000000FFF80000000003FFFFC00000;
                char[32]   <=128'h00000001FFE00000000007FFFFC00000;
                char[33]   <=128'h00000007FFC00000000007FFFFC00000;
                char[34]   <=128'h0000000FFF800000000007FFFFC00000;
                char[35]   <=128'h0000001FFF000000000003FFFF800000;
                char[36]   <=128'h0000003FFE000000000003FFFF000000;
                char[37]   <=128'h000000FFFC000000000000FFFC000000;
                char[38]   <=128'h000001FFF80000000000000000000000;
                char[39]   <=128'h000003FFF80000000000000000000000;
                char[40]   <=128'h000003FFF00000000000000000000000;
                char[41]   <=128'h000007FFF00000000000000000000000;
                char[42]   <=128'h00000FFFE00000000000000000000000;
                char[43]   <=128'h00001FFFE00000000000000000000000;
                char[44]   <=128'h00001FFFC00000000000000000000000;
                char[45]   <=128'h00003FFFC00000000000000000000000;
                char[46]   <=128'h00007FFFC00000000000000000000000;
                char[47]   <=128'h00007FFF800000000000000000000000;
                char[48]   <=128'h0000FFFF800000000000000000000000;
                char[49]   <=128'h0000FFFF800000000000000000000000;
                char[50]   <=128'h0001FFFF000000000000000000000000;
                char[51]   <=128'h0001FFFF000000000000000000000000;
                char[52]   <=128'h0001FFFF000000000000000000000000;
                char[53]   <=128'h0003FFFF000000000000000000000000;
                char[54]   <=128'h0003FFFF0000007FFFFFF80000000000;
                char[55]   <=128'h0003FFFF00000FFFFFFFFFE000000000;
                char[56]   <=128'h0007FFFF0000FFFFFFFFFFFC00000000;
                char[57]   <=128'h0007FFFE0007FFFFFFFFFFFF80000000;
                char[58]   <=128'h0007FFFE001FFFFFFFFFFFFFF0000000;
                char[59]   <=128'h0007FFFE007FFF800001FFFFF8000000;
                char[60]   <=128'h0007FFFE01FFF80000003FFFFE000000;
                char[61]   <=128'h000FFFFE07FF8000000007FFFF800000;
                char[62]   <=128'h000FFFFE0FFE0000000001FFFFC00000;
                char[63]   <=128'h000FFFFE3FF000000000007FFFE00000;
                char[64]   <=128'h000FFFFE7FC000000000003FFFF00000;
                char[65]   <=128'h000FFFFEFF8000000000000FFFF80000;
                char[66]   <=128'h000FFFFFFE00000000000007FFFC0000;
                char[67]   <=128'h000FFFFFFC00000000000003FFFE0000;
                char[68]   <=128'h000FFFFFF800000000000003FFFE0000;
                char[69]   <=128'h000FFFFFE000000000000001FFFF0000;
                char[70]   <=128'h000FFFFFC000000000000000FFFF8000;
                char[71]   <=128'h000FFFFF8000000000000000FFFF8000;
                char[72]   <=128'h000FFFFF00000000000000007FFFC000;
                char[73]   <=128'h000FFFFE00000000000000007FFFC000;
                char[74]   <=128'h000FFFFE00000000000000007FFFC000;
                char[75]   <=128'h000FFFFE00000000000000003FFFE000;
                char[76]   <=128'h0007FFFE00000000000000003FFFE000;
                char[77]   <=128'h0007FFFE00000000000000003FFFE000;
                char[78]   <=128'h0007FFFE00000000000000003FFFE000;
                char[79]   <=128'h0007FFFE00000000000000003FFFE000;
                char[80]   <=128'h0007FFFF00000000000000003FFFE000;
                char[81]   <=128'h0003FFFF00000000000000003FFFE000;
                char[82]   <=128'h0003FFFF00000000000000003FFFE000;
                char[83]   <=128'h0003FFFF00000000000000003FFFE000;
                char[84]   <=128'h0001FFFF80000000000000003FFFE000;
                char[85]   <=128'h0001FFFF80000000000000003FFFC000;
                char[86]   <=128'h0000FFFF80000000000000007FFFC000;
                char[87]   <=128'h0000FFFFC0000000000000007FFFC000;
                char[88]   <=128'h00007FFFC0000000000000007FFF8000;
                char[89]   <=128'h00007FFFE0000000000000007FFF8000;
                char[90]   <=128'h00003FFFE0000000000000007FFF8000;
                char[91]   <=128'h00001FFFF000000000000000FFFF0000;
                char[92]   <=128'h00001FFFF800000000000000FFFE0000;
                char[93]   <=128'h00000FFFFC00000000000001FFFE0000;
                char[94]   <=128'h000007FFFC00000000000001FFFC0000;
                char[95]   <=128'h000003FFFE00000000000003FFF80000;
                char[96]   <=128'h000001FFFF80000000000003FFF00000;
                char[97]   <=128'h000000FFFFC0000000000007FFE00000;
                char[98]   <=128'h0000003FFFE000000000000FFFC00000;
                char[99]   <=128'h0000001FFFF800000000001FFF000000;   
                char[100]  <=128'h00000007FFFC00000000007FFE000000; 
                char[101]  <=128'h00000003FFFF0000000001FFF8000000; 
                char[102]  <=128'h00000000FFFFE000000007FFE0000000; 
                char[103]  <=128'h000000003FFFF80000001FFF80000000; 
                char[104]  <=128'h0000000007FFFF800001FFFC00000000; 
                char[105]  <=128'h0000000000FFFFFFFFFFFFE000000000; 
                char[106]  <=128'h00000000000FFFFFFFFFFF0000000000; 
                char[107]  <=128'h000000000000FFFFFFFFE00000000000; 
                char[108]  <=128'h00000000000000FFFFF8000000000000; 
                char[109]  <=128'h00000000000000000000000000000000; 
                char[110]  <=128'h00000000000000000000000000000000; 
                char[111]  <=128'h00000000000000000000000000000000; 
                char[112]  <=128'h00000000000000000000000000000000; 
                char[113]  <=128'h00000000000000000000000000000000; 
                char[114]  <=128'h00000000000000000000000000000000; 
                char[115]  <=128'h00000000000000000000000000000000; 
                char[116]  <=128'h00000000000000000000000000000000; 
                char[117]  <=128'h00000000000000000000000000000000; 
                char[118]  <=128'h00000000000000000000000000000000; 
                char[119]  <=128'h00000000000000000000000000000000; 
                char[120]  <=128'h00000000000000000000000000000000; 
                char[121]  <=128'h00000000000000000000000000000000; 
                char[122]  <=128'h00000000000000000000000000000000; 
                char[123]  <=128'h00000000000000000000000000000000; 
                char[124]  <=128'h00000000000000000000000000000000; 
                char[125]  <=128'h00000000000000000000000000000000; 
                char[126]  <=128'h00000000000000000000000000000000; 
                char[127]  <=128'h00000000000000000000000000000000;
            end  
            4'd7:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000000000000000000;
                char[22]   <=128'h000001FFFFFFFFFFFFFFFFFFFFFF8000;
                char[23]   <=128'h000001FFFFFFFFFFFFFFFFFFFFFF8000;
                char[24]   <=128'h000003FFFFFFFFFFFFFFFFFFFFFF8000;
                char[25]   <=128'h000003FFFFFFFFFFFFFFFFFFFFFF8000;
                char[26]   <=128'h000003FFFFFFFFFFFFFFFFFFFFFF0000;
                char[27]   <=128'h000007FFFFFFFFFFFFFFFFFFFFFE0000;
                char[28]   <=128'h000007FFFFFFFFFFFFFFFFFFFFFC0000;
                char[29]   <=128'h000007FFFFFFFFFFFFFFFFFFFFF80000;
                char[30]   <=128'h00000FFFFF800000000000003FF00000;
                char[31]   <=128'h00000FFFF8000000000000007FC00000;
                char[32]   <=128'h00000FFFC000000000000000FF800000;
                char[33]   <=128'h00001FFF0000000000000001FF000000;
                char[34]   <=128'h00001FFC0000000000000003FE000000;
                char[35]   <=128'h00001FF00000000000000007FC000000;
                char[36]   <=128'h00003FE0000000000000000FF8000000;
                char[37]   <=128'h00003FC0000000000000001FF0000000;
                char[38]   <=128'h00003F80000000000000003FE0000000;
                char[39]   <=128'h00007F80000000000000007FC0000000;
                char[40]   <=128'h00007F0000000000000000FF00000000;
                char[41]   <=128'h00007E0000000000000001FE00000000;
                char[42]   <=128'h0000FE0000000000000007FC00000000;
                char[43]   <=128'h0000FC000000000000000FF800000000;
                char[44]   <=128'h000000000000000000001FF000000000;
                char[45]   <=128'h000000000000000000003FE000000000;
                char[46]   <=128'h000000000000000000007FE000000000;
                char[47]   <=128'h00000000000000000000FFC000000000;
                char[48]   <=128'h00000000000000000001FF8000000000;
                char[49]   <=128'h00000000000000000003FF0000000000;
                char[50]   <=128'h00000000000000000007FE0000000000;
                char[51]   <=128'h0000000000000000000FFC0000000000;
                char[52]   <=128'h0000000000000000001FF80000000000;
                char[53]   <=128'h0000000000000000003FF00000000000;
                char[54]   <=128'h0000000000000000007FE00000000000;
                char[55]   <=128'h000000000000000000FFC00000000000;
                char[56]   <=128'h000000000000000001FFC00000000000;
                char[57]   <=128'h000000000000000003FF800000000000;
                char[58]   <=128'h000000000000000007FF000000000000;
                char[59]   <=128'h00000000000000000FFE000000000000;
                char[60]   <=128'h00000000000000001FFE000000000000;
                char[61]   <=128'h00000000000000003FFC000000000000;
                char[62]   <=128'h00000000000000007FF8000000000000;
                char[63]   <=128'h00000000000000007FF0000000000000;
                char[64]   <=128'h0000000000000000FFF0000000000000;
                char[65]   <=128'h0000000000000001FFE0000000000000;
                char[66]   <=128'h0000000000000003FFC0000000000000;
                char[67]   <=128'h0000000000000007FFC0000000000000;
                char[68]   <=128'h000000000000000FFF80000000000000;
                char[69]   <=128'h000000000000001FFF80000000000000;
                char[70]   <=128'h000000000000001FFF00000000000000;
                char[71]   <=128'h000000000000003FFF00000000000000;
                char[72]   <=128'h000000000000007FFE00000000000000;
                char[73]   <=128'h00000000000000FFFE00000000000000;
                char[74]   <=128'h00000000000001FFFC00000000000000;
                char[75]   <=128'h00000000000001FFFC00000000000000;
                char[76]   <=128'h00000000000003FFF800000000000000;
                char[77]   <=128'h00000000000007FFF800000000000000;
                char[78]   <=128'h00000000000007FFF800000000000000;
                char[79]   <=128'h0000000000000FFFF000000000000000;
                char[80]   <=128'h0000000000000FFFF000000000000000;
                char[81]   <=128'h0000000000001FFFF000000000000000;
                char[82]   <=128'h0000000000001FFFF000000000000000;
                char[83]   <=128'h0000000000003FFFE000000000000000;
                char[84]   <=128'h0000000000003FFFE000000000000000;
                char[85]   <=128'h0000000000007FFFE000000000000000;
                char[86]   <=128'h0000000000007FFFE000000000000000;
                char[87]   <=128'h000000000000FFFFE000000000000000;
                char[88]   <=128'h000000000000FFFFE000000000000000;
                char[89]   <=128'h000000000001FFFFE000000000000000;
                char[90]   <=128'h000000000001FFFFE000000000000000;
                char[91]   <=128'h000000000001FFFFF000000000000000;
                char[92]   <=128'h000000000003FFFFF000000000000000;
                char[93]   <=128'h000000000003FFFFF000000000000000;
                char[94]   <=128'h000000000003FFFFF000000000000000;
                char[95]   <=128'h000000000003FFFFF000000000000000;
                char[96]   <=128'h000000000007FFFFF000000000000000;
                char[97]   <=128'h000000000007FFFFF000000000000000;
                char[98]   <=128'h000000000007FFFFF000000000000000;
                char[99]   <=128'h000000000007FFFFF000000000000000;  
                char[100]  <=128'h000000000007FFFFF000000000000000;
                char[101]  <=128'h000000000007FFFFF000000000000000;
                char[102]  <=128'h000000000007FFFFF000000000000000;
                char[103]  <=128'h000000000007FFFFF000000000000000;
                char[104]  <=128'h000000000003FFFFF000000000000000;
                char[105]  <=128'h000000000003FFFFE000000000000000;
                char[106]  <=128'h000000000001FFFFE000000000000000;
                char[107]  <=128'h0000000000007FFFC000000000000000;
                char[108]  <=128'h0000000000000FFE0000000000000000;
                char[109]  <=128'h00000000000000000000000000000000;
                char[110]  <=128'h00000000000000000000000000000000;
                char[111]  <=128'h00000000000000000000000000000000;
                char[112]  <=128'h00000000000000000000000000000000;
                char[113]  <=128'h00000000000000000000000000000000;
                char[114]  <=128'h00000000000000000000000000000000;
                char[115]  <=128'h00000000000000000000000000000000;
                char[116]  <=128'h00000000000000000000000000000000;
                char[117]  <=128'h00000000000000000000000000000000;
                char[118]  <=128'h00000000000000000000000000000000;
                char[119]  <=128'h00000000000000000000000000000000;
                char[120]  <=128'h00000000000000000000000000000000;
                char[121]  <=128'h00000000000000000000000000000000;
                char[122]  <=128'h00000000000000000000000000000000;
                char[123]  <=128'h00000000000000000000000000000000;
                char[124]  <=128'h00000000000000000000000000000000;
                char[125]  <=128'h00000000000000000000000000000000;
                char[126]  <=128'h00000000000000000000000000000000;
                char[127]  <=128'h00000000000000000000000000000000; 
            end
            4'd8:
            begin
                char[0]    <=128'h00000000000000000000000000000000;
                char[1]    <=128'h00000000000000000000000000000000;
                char[2]    <=128'h00000000000000000000000000000000;
                char[3]    <=128'h00000000000000000000000000000000;
                char[4]    <=128'h00000000000000000000000000000000;
                char[5]    <=128'h00000000000000000000000000000000;
                char[6]    <=128'h00000000000000000000000000000000;
                char[7]    <=128'h00000000000000000000000000000000;
                char[8]    <=128'h00000000000000000000000000000000;
                char[9]    <=128'h00000000000000000000000000000000;
                char[10]   <=128'h00000000000000000000000000000000;
                char[11]   <=128'h00000000000000000000000000000000;
                char[12]   <=128'h00000000000000000000000000000000;
                char[13]   <=128'h00000000000000000000000000000000;
                char[14]   <=128'h00000000000000000000000000000000;
                char[15]   <=128'h00000000000000000000000000000000;
                char[16]   <=128'h00000000000000000000000000000000;
                char[17]   <=128'h00000000000000000000000000000000;
                char[18]   <=128'h00000000000000000000000000000000;
                char[19]   <=128'h00000000000000000000000000000000;
                char[20]   <=128'h00000000000000000000000000000000;
                char[21]   <=128'h00000000000000000000000000000000;
                char[22]   <=128'h000000000001FFFFFFFF000000000000;
                char[23]   <=128'h00000000007FFFFFFFFFFC0000000000;
                char[24]   <=128'h000000000FFFFFFFFFFFFFC000000000;
                char[25]   <=128'h000000007FFFF800003FFFF800000000;
                char[26]   <=128'h00000003FFFC00000000FFFF00000000;
                char[27]   <=128'h0000000FFFE0000000001FFFC0000000;
                char[28]   <=128'h0000003FFF000000000003FFF0000000;
                char[29]   <=128'h000000FFFC000000000000FFFC000000;
                char[30]   <=128'h000001FFF00000000000007FFE000000;
                char[31]   <=128'h000007FFE00000000000001FFF800000;
                char[32]   <=128'h00000FFFC00000000000000FFFC00000;
                char[33]   <=128'h00001FFF0000000000000007FFE00000;
                char[34]   <=128'h00003FFF0000000000000003FFF00000;
                char[35]   <=128'h00007FFE0000000000000001FFF80000;
                char[36]   <=128'h00007FFC0000000000000001FFF80000;
                char[37]   <=128'h0000FFFC0000000000000000FFFC0000;
                char[38]   <=128'h0000FFF80000000000000000FFFC0000;
                char[39]   <=128'h0001FFF800000000000000007FFE0000;
                char[40]   <=128'h0001FFF800000000000000007FFE0000;
                char[41]   <=128'h0001FFF800000000000000007FFE0000;
                char[42]   <=128'h0001FFF800000000000000007FFE0000;
                char[43]   <=128'h0001FFFC00000000000000007FFE0000;
                char[44]   <=128'h0001FFFE00000000000000007FFE0000;
                char[45]   <=128'h0000FFFE00000000000000007FFC0000;
                char[46]   <=128'h0000FFFF8000000000000000FFFC0000;
                char[47]   <=128'h0000FFFFC000000000000000FFF80000;
                char[48]   <=128'h00007FFFE000000000000001FFF80000;
                char[49]   <=128'h00003FFFF800000000000001FFF00000;
                char[50]   <=128'h00001FFFFE00000000000003FFE00000;
                char[51]   <=128'h00000FFFFF80000000000007FFC00000;
                char[52]   <=128'h000007FFFFE000000000000FFF800000;
                char[53]   <=128'h000003FFFFFC00000000003FFE000000;
                char[54]   <=128'h000000FFFFFF80000000007FFC000000;
                char[55]   <=128'h0000007FFFFFF000000001FFF0000000;
                char[56]   <=128'h0000001FFFFFFE00000007FFC0000000;
                char[57]   <=128'h00000007FFFFFFE000001FFF00000000;
                char[58]   <=128'h00000001FFFFFFFE0000FFF800000000;
                char[59]   <=128'h000000003FFFFFFFF007FFC000000000;
                char[60]   <=128'h0000000007FFFFFFFFFFFE0000000000;
                char[61]   <=128'h0000000000FFFFFFFFFFF00000000000;
                char[62]   <=128'h00000000000FFFFFFFFF000000000000;
                char[63]   <=128'h00000000007FFFFFFFFFE00000000000;
                char[64]   <=128'h0000000007FFFFFFFFFFFC0000000000;
                char[65]   <=128'h000000001FFE01FFFFFFFF8000000000;
                char[66]   <=128'h00000000FFF8001FFFFFFFF000000000;
                char[67]   <=128'h00000003FFC00001FFFFFFFC00000000;
                char[68]   <=128'h0000001FFF0000001FFFFFFF00000000;
                char[69]   <=128'h0000007FFC00000003FFFFFFC0000000;
                char[70]   <=128'h000001FFF8000000007FFFFFF0000000;
                char[71]   <=128'h000003FFE0000000000FFFFFFC000000;
                char[72]   <=128'h00000FFFC00000000001FFFFFF000000;
                char[73]   <=128'h00001FFF8000000000003FFFFF800000;
                char[74]   <=128'h00003FFF0000000000000FFFFFC00000;
                char[75]   <=128'h0000FFFC00000000000003FFFFE00000;
                char[76]   <=128'h0001FFFC00000000000000FFFFF00000;
                char[77]   <=128'h0001FFF8000000000000003FFFF80000;
                char[78]   <=128'h0003FFF0000000000000001FFFFC0000;
                char[79]   <=128'h0007FFE00000000000000007FFFE0000;
                char[80]   <=128'h0007FFE00000000000000003FFFE0000;
                char[81]   <=128'h000FFFC00000000000000001FFFF0000;
                char[82]   <=128'h000FFFC00000000000000000FFFF0000;
                char[83]   <=128'h000FFFC000000000000000007FFF8000;
                char[84]   <=128'h001FFF8000000000000000007FFF8000;
                char[85]   <=128'h001FFF8000000000000000003FFF8000;
                char[86]   <=128'h001FFF8000000000000000003FFF8000;
                char[87]   <=128'h001FFF8000000000000000003FFF8000;
                char[88]   <=128'h001FFF8000000000000000003FFF8000;
                char[89]   <=128'h001FFF8000000000000000003FFF8000;
                char[90]   <=128'h001FFF8000000000000000003FFF0000;
                char[91]   <=128'h000FFFC000000000000000007FFF0000;
                char[92]   <=128'h000FFFC000000000000000007FFE0000;
                char[93]   <=128'h0007FFE000000000000000007FFE0000;
                char[94]   <=128'h0003FFE00000000000000000FFFC0000;
                char[95]   <=128'h0001FFF00000000000000001FFF80000;
                char[96]   <=128'h0000FFF80000000000000001FFF00000;
                char[97]   <=128'h00007FFC0000000000000003FFE00000;
                char[98]   <=128'h00003FFF000000000000000FFFC00000;
                char[99]   <=128'h00000FFFC00000000000001FFF000000;   
                char[100]  <=128'h000003FFF00000000000007FFE000000; 
                char[101]  <=128'h000000FFFC000000000000FFF8000000; 
                char[102]  <=128'h0000003FFF800000000007FFE0000000; 
                char[103]  <=128'h0000000FFFF0000000003FFF80000000; 
                char[104]  <=128'h00000001FFFF80000007FFFC00000000; 
                char[105]  <=128'h000000003FFFFFFFFFFFFFE000000000; 
                char[106]  <=128'h0000000003FFFFFFFFFFFE0000000000; 
                char[107]  <=128'h00000000001FFFFFFFFFC00000000000; 
                char[108]  <=128'h0000000000001FFFFFC0000000000000; 
                char[109]  <=128'h00000000000000000000000000000000; 
                char[110]  <=128'h00000000000000000000000000000000; 
                char[111]  <=128'h00000000000000000000000000000000; 
                char[112]  <=128'h00000000000000000000000000000000; 
                char[113]  <=128'h00000000000000000000000000000000; 
                char[114]  <=128'h00000000000000000000000000000000; 
                char[115]  <=128'h00000000000000000000000000000000; 
                char[116]  <=128'h00000000000000000000000000000000; 
                char[117]  <=128'h00000000000000000000000000000000; 
                char[118]  <=128'h00000000000000000000000000000000; 
                char[119]  <=128'h00000000000000000000000000000000; 
                char[120]  <=128'h00000000000000000000000000000000; 
                char[121]  <=128'h00000000000000000000000000000000; 
                char[122]  <=128'h00000000000000000000000000000000; 
                char[123]  <=128'h00000000000000000000000000000000; 
                char[124]  <=128'h00000000000000000000000000000000; 
                char[125]  <=128'h00000000000000000000000000000000; 
                char[126]  <=128'h00000000000000000000000000000000; 
                char[127]  <=128'h00000000000000000000000000000000;  
            end
            4'd9:
        begin
            char[0]    <=128'h00000000000000000000000000000000;
            char[1]    <=128'h00000000000000000000000000000000;
            char[2]    <=128'h00000000000000000000000000000000;
            char[3]    <=128'h00000000000000000000000000000000;
            char[4]    <=128'h00000000000000000000000000000000;
            char[5]    <=128'h00000000000000000000000000000000;
            char[6]    <=128'h00000000000000000000000000000000;
            char[7]    <=128'h00000000000000000000000000000000;
            char[8]    <=128'h00000000000000000000000000000000;
            char[9]    <=128'h00000000000000000000000000000000;
            char[10]   <=128'h00000000000000000000000000000000;
            char[11]   <=128'h00000000000000000000000000000000;
            char[12]   <=128'h00000000000000000000000000000000;
            char[13]   <=128'h00000000000000000000000000000000;
            char[14]   <=128'h00000000000000000000000000000000;
            char[15]   <=128'h00000000000000000000000000000000;
            char[16]   <=128'h00000000000000000000000000000000;
            char[17]   <=128'h00000000000000000000000000000000;
            char[18]   <=128'h00000000000000000000000000000000;
            char[19]   <=128'h00000000000000000000000000000000;
            char[20]   <=128'h00000000000000000000000000000000;
            char[21]   <=128'h00000000000000000000000000000000;
            char[22]   <=128'h000000000007FFFFFFF0000000000000;
            char[23]   <=128'h0000000000FFFFFFFFFF800000000000;
            char[24]   <=128'h000000000FFFFFFFFFFFF80000000000;
            char[25]   <=128'h000000007FFFF00003FFFF0000000000;
            char[26]   <=128'h00000003FFFE0000001FFFE000000000;
            char[27]   <=128'h0000000FFFF000000001FFF800000000;
            char[28]   <=128'h0000003FFF80000000007FFE00000000;
            char[29]   <=128'h000000FFFE00000000001FFF80000000;
            char[30]   <=128'h000003FFFC000000000007FFE0000000;
            char[31]   <=128'h000007FFF0000000000003FFF0000000;
            char[32]   <=128'h00000FFFE0000000000001FFF8000000;
            char[33]   <=128'h00001FFFC0000000000000FFFE000000;
            char[34]   <=128'h00003FFF800000000000007FFF000000;
            char[35]   <=128'h00007FFF000000000000003FFF800000;
            char[36]   <=128'h0000FFFF000000000000001FFFC00000;
            char[37]   <=128'h0001FFFE000000000000001FFFC00000;
            char[38]   <=128'h0003FFFC000000000000000FFFE00000;
            char[39]   <=128'h0003FFFC000000000000000FFFF00000;
            char[40]   <=128'h0007FFFC0000000000000007FFF80000;
            char[41]   <=128'h0007FFF80000000000000007FFF80000;
            char[42]   <=128'h000FFFF80000000000000003FFFC0000;
            char[43]   <=128'h000FFFF80000000000000003FFFC0000;
            char[44]   <=128'h000FFFF00000000000000003FFFE0000;
            char[45]   <=128'h001FFFF00000000000000003FFFE0000;
            char[46]   <=128'h001FFFF00000000000000001FFFF0000;
            char[47]   <=128'h001FFFF00000000000000001FFFF0000;
            char[48]   <=128'h001FFFF00000000000000001FFFF0000;
            char[49]   <=128'h001FFFF00000000000000001FFFF8000;
            char[50]   <=128'h001FFFF00000000000000001FFFF8000;
            char[51]   <=128'h001FFFF00000000000000001FFFF8000;
            char[52]   <=128'h001FFFF00000000000000001FFFF8000;
            char[53]   <=128'h001FFFF00000000000000001FFFF8000;
            char[54]   <=128'h001FFFF80000000000000003FFFFC000;
            char[55]   <=128'h000FFFF80000000000000003FFFFC000;
            char[56]   <=128'h000FFFF80000000000000007FFFFC000;
            char[57]   <=128'h000FFFFC000000000000000FFFFFC000;
            char[58]   <=128'h0007FFFC000000000000000FFFFFC000;
            char[59]   <=128'h0007FFFE000000000000001FFFFFC000;
            char[60]   <=128'h0007FFFE000000000000007FFFFFC000;
            char[61]   <=128'h0003FFFF00000000000000FFFFFFC000;
            char[62]   <=128'h0001FFFF80000000000001FFFFFFC000;
            char[63]   <=128'h0001FFFFC0000000000003FDFFFFC000;
            char[64]   <=128'h0000FFFFE000000000000FF9FFFFC000;
            char[65]   <=128'h00007FFFF000000000003FE1FFFFC000;
            char[66]   <=128'h00003FFFFC0000000000FFC1FFFFC000;
            char[67]   <=128'h00001FFFFE0000000003FF83FFFFC000;
            char[68]   <=128'h000007FFFFC00000000FFE03FFFF8000;
            char[69]   <=128'h000001FFFFF00000007FF803FFFF8000;
            char[70]   <=128'h0000007FFFFF000007FFE003FFFF8000;
            char[71]   <=128'h0000001FFFFFFFFFFFFF8003FFFF8000;
            char[72]   <=128'h00000003FFFFFFFFFFFE0003FFFF8000;
            char[73]   <=128'h000000007FFFFFFFFFF00007FFFF0000;
            char[74]   <=128'h0000000007FFFFFFFE000007FFFF0000;
            char[75]   <=128'h00000000000FFFFF80000007FFFF0000;
            char[76]   <=128'h000000000000000000000007FFFE0000;
            char[77]   <=128'h00000000000000000000000FFFFE0000;
            char[78]   <=128'h00000000000000000000000FFFFC0000;
            char[79]   <=128'h00000000000000000000000FFFFC0000;
            char[80]   <=128'h00000000000000000000001FFFF80000;
            char[81]   <=128'h00000000000000000000001FFFF80000;
            char[82]   <=128'h00000000000000000000001FFFF00000;
            char[83]   <=128'h00000000000000000000003FFFF00000;
            char[84]   <=128'h00000000000000000000003FFFE00000;
            char[85]   <=128'h00000000000000000000007FFFE00000;
            char[86]   <=128'h00000000000000000000007FFFC00000;
            char[87]   <=128'h0000000000000000000000FFFF800000;
            char[88]   <=128'h0000000000000000000000FFFF000000;
            char[89]   <=128'h0000000000000000000001FFFE000000;
            char[90]   <=128'h0000000000000000000003FFFE000000;
            char[91]   <=128'h0000000000000000000003FFFC000000;
            char[92]   <=128'h0000003FF0000000000007FFF8000000;
            char[93]   <=128'h000001FFFC00000000000FFFF0000000;
            char[94]   <=128'h000003FFFE00000000001FFFC0000000;
            char[95]   <=128'h000007FFFF00000000003FFF80000000;
            char[96]   <=128'h00000FFFFF00000000007FFF00000000;
            char[97]   <=128'h00000FFFFF8000000000FFFE00000000;
            char[98]   <=128'h00000FFFFF8000000003FFF800000000;
            char[99]   <=128'h00000FFFFF8000000007FFF000000000;   
            char[100]  <=128'h000007FFFF800000001FFFC000000000; 
            char[101]  <=128'h000007FFFF800000007FFF0000000000; 
            char[102]  <=128'h000003FFFFC0000001FFFC0000000000; 
            char[103]  <=128'h000000FFFFE000000FFFF00000000000; 
            char[104]  <=128'h0000003FFFF00000FFFF800000000000; 
            char[105]  <=128'h0000000FFFFFFFFFFFFC000000000000; 
            char[106]  <=128'h00000001FFFFFFFFFFC0000000000000; 
            char[107]  <=128'h000000001FFFFFFFFC00000000000000; 
            char[108]  <=128'h00000000003FFFFE0000000000000000; 
            char[109]  <=128'h00000000000000000000000000000000; 
            char[110]  <=128'h00000000000000000000000000000000; 
            char[111]  <=128'h00000000000000000000000000000000; 
            char[112]  <=128'h00000000000000000000000000000000; 
            char[113]  <=128'h00000000000000000000000000000000; 
            char[114]  <=128'h00000000000000000000000000000000; 
            char[115]  <=128'h00000000000000000000000000000000; 
            char[116]  <=128'h00000000000000000000000000000000; 
            char[117]  <=128'h00000000000000000000000000000000; 
            char[118]  <=128'h00000000000000000000000000000000; 
            char[119]  <=128'h00000000000000000000000000000000; 
            char[120]  <=128'h00000000000000000000000000000000; 
            char[121]  <=128'h00000000000000000000000000000000; 
            char[122]  <=128'h00000000000000000000000000000000; 
            char[123]  <=128'h00000000000000000000000000000000; 
            char[124]  <=128'h00000000000000000000000000000000; 
            char[125]  <=128'h00000000000000000000000000000000; 
            char[126]  <=128'h00000000000000000000000000000000; 
            char[127]  <=128'h00000000000000000000000000000000;  
        end
            4'd10:
        begin
            char[0]    <={32'h00000000,96'h0};
            char[1]    <={32'h00000000,96'h0};
            char[2]    <={32'h00000000,96'h0};
            char[3]    <={32'h00000000,96'h0};
            char[4]    <={32'h00000000,96'h0};
            char[5]    <={32'h00000000,96'h0};
            char[6]    <={32'h00000000,96'h0};
            char[7]    <={32'h00000000,96'h0};
            char[8]    <={32'h00000000,96'h0};
            char[9]    <={32'h00000000,96'h0};
            char[10]   <={32'h00000000,96'h0};
            char[11]   <={32'h00000000,96'h0};
            char[12]   <={32'h00000000,96'h0};
            char[13]   <={32'h00000000,96'h0};
            char[14]   <={32'h00000000,96'h0};
            char[15]   <={32'h00000000,96'h0};
            char[16]   <={32'h00000000,96'h0};
            char[17]   <={32'h00000000,96'h0};
            char[18]   <={32'h00000000,96'h0};
            char[19]   <={32'h00000000,96'h0};
            char[20]   <={32'h00000000,96'h0};
            char[21]   <={32'h00000000,96'h0};
            char[22]   <={32'h00000000,96'h0};
            char[23]   <={32'h00000000,96'h0};
            char[24]   <={32'h00000000,96'h0};
            char[25]   <={32'h00000000,96'h0};
            char[26]   <={32'h00000000,96'h0};
            char[27]   <={32'h00000000,96'h0};
            char[28]   <={32'h00000000,96'h0};
            char[29]   <={32'h00000000,96'h0};
            char[30]   <={32'h00000000,96'h0};
            char[31]   <={32'h00000000,96'h0};
            char[32]   <={32'h00000000,96'h0};
            char[33]   <={32'h00000000,96'h0};
            char[34]   <={32'h00000000,96'h0};
            char[35]   <={32'h00000000,96'h0};
            char[36]   <={32'h00000000,96'h0};
            char[37]   <={32'h00000000,96'h0};
            char[38]   <={32'h00000000,96'h0};
            char[39]   <={32'h00000000,96'h0};
            char[40]   <={32'h00000000,96'h0};
            char[41]   <={32'h0001E000,96'h0};
            char[42]   <={32'h0003F000,96'h0};
            char[43]   <={32'h0007F000,96'h0};
            char[44]   <={32'h0007F800,96'h0};
            char[45]   <={32'h000FF800,96'h0};
            char[46]   <={32'h000FF800,96'h0};
            char[47]   <={32'h000FF800,96'h0};
            char[48]   <={32'h000FF800,96'h0};
            char[49]   <={32'h000FF800,96'h0};
            char[50]   <={32'h000FF800,96'h0};
            char[51]   <={32'h000FF800,96'h0};
            char[52]   <={32'h000FF800,96'h0};
            char[53]   <={32'h0007F800,96'h0};
            char[54]   <={32'h0007F000,96'h0};
            char[55]   <={32'h0007F000,96'h0};
            char[56]   <={32'h0003E000,96'h0};
            char[57]   <={32'h0001C000,96'h0};
            char[58]   <={32'h00000000,96'h0};
            char[59]   <={32'h00000000,96'h0};
            char[60]   <={32'h00000000,96'h0};
            char[61]   <={32'h00000000,96'h0};
            char[62]   <={32'h00000000,96'h0};
            char[63]   <={32'h00000000,96'h0};
            char[64]   <={32'h00000000,96'h0};
            char[65]   <={32'h00000000,96'h0};
            char[66]   <={32'h00000000,96'h0};
            char[67]   <={32'h00000000,96'h0};
            char[68]   <={32'h00000000,96'h0};
            char[69]   <={32'h00000000,96'h0};
            char[70]   <={32'h00008000,96'h0};
            char[71]   <={32'h0003E000,96'h0};
            char[72]   <={32'h0007F000,96'h0};
            char[73]   <={32'h0007F000,96'h0};
            char[74]   <={32'h0007F000,96'h0};
            char[75]   <={32'h000FF800,96'h0};
            char[76]   <={32'h000FF800,96'h0};
            char[77]   <={32'h000FF800,96'h0};
            char[78]   <={32'h000FF800,96'h0};
            char[79]   <={32'h000FF800,96'h0};
            char[80]   <={32'h000FF800,96'h0};
            char[81]   <={32'h000FF800,96'h0};
            char[82]   <={32'h000FF800,96'h0};
            char[83]   <={32'h0007F000,96'h0};
            char[84]   <={32'h0007F000,96'h0};
            char[85]   <={32'h0003E000,96'h0};
            char[86]   <={32'h0003E000,96'h0};
            char[87]   <={32'h00008000,96'h0};
            char[88]   <={32'h00000000,96'h0};
            char[89]   <={32'h00000000,96'h0};
            char[90]   <={32'h00000000,96'h0};
            char[91]   <={32'h00000000,96'h0};
            char[92]   <={32'h00000000,96'h0};
            char[93]   <={32'h00000000,96'h0};
            char[94]   <={32'h00000000,96'h0};
            char[95]   <={32'h00000000,96'h0};
            char[96]   <={32'h00000000,96'h0};
            char[97]   <={32'h00000000,96'h0};
            char[98]   <={32'h00000000,96'h0};
            char[99]   <={32'h00000000,96'h0};   
            char[100]  <={32'h00000000,96'h0}; 
            char[101]  <={32'h00000000,96'h0}; 
            char[102]  <={32'h00000000,96'h0}; 
            char[103]  <={32'h00000000,96'h0}; 
            char[104]  <={32'h00000000,96'h0}; 
            char[105]  <={32'h00000000,96'h0}; 
            char[106]  <={32'h00000000,96'h0}; 
            char[107]  <={32'h00000000,96'h0}; 
            char[108]  <={32'h00000000,96'h0}; 
            char[109]  <={32'h00000000,96'h0}; 
            char[110]  <={32'h00000000,96'h0}; 
            char[111]  <={32'h00000000,96'h0}; 
            char[112]  <={32'h00000000,96'h0}; 
            char[113]  <={32'h00000000,96'h0}; 
            char[114]  <={32'h00000000,96'h0}; 
            char[115]  <={32'h00000000,96'h0}; 
            char[116]  <={32'h00000000,96'h0}; 
            char[117]  <={32'h00000000,96'h0}; 
            char[118]  <={32'h00000000,96'h0}; 
            char[119]  <={32'h00000000,96'h0}; 
            char[120]  <={32'h00000000,96'h0}; 
            char[121]  <={32'h00000000,96'h0}; 
            char[122]  <={32'h00000000,96'h0}; 
            char[123]  <={32'h00000000,96'h0}; 
            char[124]  <={32'h00000000,96'h0}; 
            char[125]  <={32'h00000000,96'h0}; 
            char[126]  <={32'h00000000,96'h0}; 
            char[127]  <={32'h00000000,96'h0};  
        end
        default:;
        endcase
end


// 当收到字符数据请求的时候，向外部输出char_data的数据。
always @(posedge clk or negedge rst_n) begin
    if (~rst_n)
        char_data <= 1'b0;
    else if(char_data_req)
        char_data <= char[char_y_loc][127-char_x_loc];
end

endmodule